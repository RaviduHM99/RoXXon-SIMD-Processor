`timescale 1ns/1ps

module Fetch_Unit #(
    parameter N = 2
)(
    input logic CLK, RSTN,

);


endmodule