`timescale 1ns/1ps

module Instruction_RF #(
    parameter N = 512
)(
    input logic CLK,

    output logic [31:0] INSTR_AXI,
    input logic [$clog2(N)-1:0] PC_AXI

);

    reg [16:0][31:0] AXI_SLAVE_REG;

    initial begin
      /* 
        ////////////////////////////////////////////////////////////////////////
        //////////////// 8x8 Matrix Multiplication Instructions ////////////////
        ////////////////////////////////////////////////////////////////////////

        AXI_SLAVE_REG[0] <= 32'b0000_00_0000_00_0_0_10_010; //LOADA Row1
        AXI_SLAVE_REG[1] <= 32'b1000000_00_0000_01_0_0_10_011; //LOADB Col1
        AXI_SLAVE_REG[2] <= 32'b1001000_01_0000_01_0_0_10_011; //LOADB Col2
        AXI_SLAVE_REG[3] <= 32'b1010000_10_0000_01_0_0_10_011; //LOADB Col3
        AXI_SLAVE_REG[4] <= 32'b1011000_11_0000_01_0_0_10_011; //LOADB Col4
        AXI_SLAVE_REG[5] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[6] <= 32'b10000000_00_0000_00_0_0_10_101; //STORE Row1 - 1/2
        AXI_SLAVE_REG[7] <= 32'b1100000_00_0000_01_0_1_10_011; //LOADB Col5
        AXI_SLAVE_REG[8] <= 32'b1101000_01_0000_01_0_0_10_011; //LOADB Col6
        AXI_SLAVE_REG[9] <= 32'b1110000_10_0000_01_0_0_10_011; //LOADB Col7
        AXI_SLAVE_REG[10] <= 32'b1111000_11_0000_01_0_0_10_011; //LOADB Col8
        AXI_SLAVE_REG[11] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[12] <= 32'b10001000_00_0000_00_0_0_10_101; //STORE Row1 - 2/2

        AXI_SLAVE_REG[13] <= 32'b0000_00_0000_00_0_0_10_010; //LOADA Row2
        AXI_SLAVE_REG[14] <= 32'b1000000_00_0000_01_0_0_10_011; //LOADB Col1
        AXI_SLAVE_REG[15] <= 32'b1001000_01_0000_01_0_0_10_011; //LOADB Col2
        AXI_SLAVE_REG[16] <= 32'b1010000_10_0000_01_0_0_10_011; //LOADB Col3
        AXI_SLAVE_REG[17] <= 32'b1011000_11_0000_01_0_0_10_011; //LOADB Col4
        AXI_SLAVE_REG[18] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[19] <= 32'b10010000_00_0000_00_0_0_10_101; //STORE Row2 - 1/2
        AXI_SLAVE_REG[20] <= 32'b1100000_00_0000_01_0_1_10_011; //LOADB Col5
        AXI_SLAVE_REG[21] <= 32'b1101000_01_0000_01_0_0_10_011; //LOADB Col6
        AXI_SLAVE_REG[22] <= 32'b1110000_10_0000_01_0_0_10_011; //LOADB Col7
        AXI_SLAVE_REG[23] <= 32'b1111000_11_0000_01_0_0_10_011; //LOADB Col8
        AXI_SLAVE_REG[24] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[25] <= 32'b10011000_00_0000_00_0_0_10_101; //STORE Row2 - 2/2

        AXI_SLAVE_REG[26] <= 32'b0000_00_0000_00_0_0_10_010; //LOADA Row3
        AXI_SLAVE_REG[27] <= 32'b1000000_00_0000_01_0_0_10_011; //LOADB Col1
        AXI_SLAVE_REG[28] <= 32'b1001000_01_0000_01_0_0_10_011; //LOADB Col2
        AXI_SLAVE_REG[29] <= 32'b1010000_10_0000_01_0_0_10_011; //LOADB Col3
        AXI_SLAVE_REG[30] <= 32'b1011000_11_0000_01_0_0_10_011; //LOADB Col4
        AXI_SLAVE_REG[31] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[32] <= 32'b10100000_00_0000_00_0_0_10_101; //STORE Row3 - 1/2
        AXI_SLAVE_REG[33] <= 32'b1100000_00_0000_01_0_1_10_011; //LOADB Col5
        AXI_SLAVE_REG[34] <= 32'b1101000_01_0000_01_0_0_10_011; //LOADB Col6
        AXI_SLAVE_REG[35] <= 32'b1110000_10_0000_01_0_0_10_011; //LOADB Col7
        AXI_SLAVE_REG[36] <= 32'b1111000_11_0000_01_0_0_10_011; //LOADB Col8
        AXI_SLAVE_REG[37] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[38] <= 32'b10101000_00_0000_00_0_0_10_101; //STORE Row3 - 2/2

        AXI_SLAVE_REG[39] <= 32'b0000_00_0000_00_0_0_10_010; //LOADA Row4
        AXI_SLAVE_REG[40] <= 32'b1000000_00_0000_01_0_0_10_011; //LOADB Col1
        AXI_SLAVE_REG[41] <= 32'b1001000_01_0000_01_0_0_10_011; //LOADB Col2
        AXI_SLAVE_REG[42] <= 32'b1010000_10_0000_01_0_0_10_011; //LOADB Col3
        AXI_SLAVE_REG[43] <= 32'b1011000_11_0000_01_0_0_10_011; //LOADB Col4
        AXI_SLAVE_REG[44] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[45] <= 32'b10110000_00_0000_00_0_0_10_101; //STORE Row4 - 1/2
        AXI_SLAVE_REG[46] <= 32'b1100000_00_0000_01_0_1_10_011; //LOADB Col5
        AXI_SLAVE_REG[47] <= 32'b1101000_01_0000_01_0_0_10_011; //LOADB Col6
        AXI_SLAVE_REG[48] <= 32'b1110000_10_0000_01_0_0_10_011; //LOADB Col7
        AXI_SLAVE_REG[49] <= 32'b1111000_11_0000_01_0_0_10_011; //LOADB Col8
        AXI_SLAVE_REG[50] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[51] <= 32'b10111000_00_0000_00_0_0_10_101; //STORE Row4 - 2/2

        AXI_SLAVE_REG[52] <= 32'b0000_00_0000_00_0_0_10_010; //LOADA Row5
        AXI_SLAVE_REG[53] <= 32'b1000000_00_0000_01_0_0_10_011; //LOADB Col1
        AXI_SLAVE_REG[54] <= 32'b1001000_01_0000_01_0_0_10_011; //LOADB Col2
        AXI_SLAVE_REG[55] <= 32'b1010000_10_0000_01_0_0_10_011; //LOADB Col3
        AXI_SLAVE_REG[56] <= 32'b1011000_11_0000_01_0_0_10_011; //LOADB Col4
        AXI_SLAVE_REG[57] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[58] <= 32'b100000_00_0000_00_0_0_10_101; //STORE Row5 - 1/2
        AXI_SLAVE_REG[59] <= 32'b1100000_00_0000_01_0_1_10_011; //LOADB Col5
        AXI_SLAVE_REG[60] <= 32'b1101000_01_0000_01_0_0_10_011; //LOADB Col6
        AXI_SLAVE_REG[61] <= 32'b1110000_10_0000_01_0_0_10_011; //LOADB Col7
        AXI_SLAVE_REG[62] <= 32'b1111000_11_0000_01_0_0_10_011; //LOADB Col8
        AXI_SLAVE_REG[63] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[64] <= 32'b100000_00_0000_00_0_0_10_101; //STORE Row5 - 2/2

        AXI_SLAVE_REG[65] <= 32'b0000_00_0000_00_0_0_10_010; //LOADA Row6
        AXI_SLAVE_REG[66] <= 32'b1000000_00_0000_01_0_0_10_011; //LOADB Col1
        AXI_SLAVE_REG[67] <= 32'b1001000_01_0000_01_0_0_10_011; //LOADB Col2
        AXI_SLAVE_REG[68] <= 32'b1010000_10_0000_01_0_0_10_011; //LOADB Col3
        AXI_SLAVE_REG[69] <= 32'b1011000_11_0000_01_0_0_10_011; //LOADB Col4
        AXI_SLAVE_REG[70] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[71] <= 32'b100000_00_0000_00_0_0_10_101; //STORE Row6 - 1/2
        AXI_SLAVE_REG[72] <= 32'b1100000_00_0000_01_0_1_10_011; //LOADB Col5
        AXI_SLAVE_REG[73] <= 32'b1101000_01_0000_01_0_0_10_011; //LOADB Col6
        AXI_SLAVE_REG[74] <= 32'b1110000_10_0000_01_0_0_10_011; //LOADB Col7
        AXI_SLAVE_REG[75] <= 32'b1111000_11_0000_01_0_0_10_011; //LOADB Col8
        AXI_SLAVE_REG[76] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[77] <= 32'b100000_00_0000_00_0_0_10_101; //STORE Row6 - 2/2

        AXI_SLAVE_REG[78] <= 32'b0000_00_0000_00_0_0_10_010; //LOADA Row7
        AXI_SLAVE_REG[79] <= 32'b1000000_00_0000_01_0_0_10_011; //LOADB Col1
        AXI_SLAVE_REG[80] <= 32'b1001000_01_0000_01_0_0_10_011; //LOADB Col2
        AXI_SLAVE_REG[81] <= 32'b1010000_10_0000_01_0_0_10_011; //LOADB Col3
        AXI_SLAVE_REG[82] <= 32'b1011000_11_0000_01_0_0_10_011; //LOADB Col4
        AXI_SLAVE_REG[83] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[84] <= 32'b100000_00_0000_00_0_0_10_101; //STORE Row7 - 1/2
        AXI_SLAVE_REG[85] <= 32'b1100000_00_0000_01_0_1_10_011; //LOADB Col5
        AXI_SLAVE_REG[86] <= 32'b1101000_01_0000_01_0_0_10_011; //LOADB Col6
        AXI_SLAVE_REG[87] <= 32'b1110000_10_0000_01_0_0_10_011; //LOADB Col7
        AXI_SLAVE_REG[88] <= 32'b1111000_11_0000_01_0_0_10_011; //LOADB Col8
        AXI_SLAVE_REG[89] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[90] <= 32'b100000_00_0000_00_0_0_10_101; //STORE Row7 - 2/2

        AXI_SLAVE_REG[91] <= 32'b0000_00_0000_00_0_0_10_010; //LOADA Row8
        AXI_SLAVE_REG[92] <= 32'b1000000_00_0000_01_0_0_10_011; //LOADB Col1
        AXI_SLAVE_REG[93] <= 32'b1001000_01_0000_01_0_0_10_011; //LOADB Col2
        AXI_SLAVE_REG[94] <= 32'b1010000_10_0000_01_0_0_10_011; //LOADB Col3
        AXI_SLAVE_REG[95] <= 32'b1011000_11_0000_01_0_0_10_011; //LOADB Col4
        AXI_SLAVE_REG[96] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[97] <= 32'b100000_00_0000_00_0_0_10_101; //STORE Row8 - 1/2
        AXI_SLAVE_REG[98] <= 32'b1100000_00_0000_01_0_1_10_011; //LOADB Col5
        AXI_SLAVE_REG[99] <= 32'b1101000_01_0000_01_0_0_10_011; //LOADB Col6
        AXI_SLAVE_REG[100] <= 32'b1110000_10_0000_01_0_0_10_011; //LOADB Col7
        AXI_SLAVE_REG[101] <= 32'b1111000_11_0000_01_0_0_10_011; //LOADB Col8
        AXI_SLAVE_REG[102] <= 32'b0000_00_0000_01_0_0_10_100; //MULTACC
        AXI_SLAVE_REG[103] <= 32'b100000_00_0000_00_0_0_10_101; //STORE Row8 - 2/2

        AXI_SLAVE_REG[104] <= 32'b0000_00_0000_00_0_0_00_110; //STOP 
*/
        ////////////////////////////////////////////////////////////////////////
        //////////////// 4x4 Matrix Multiplication Instructions ////////////////
        ////////////////////////////////////////////////////////////////////////
    
        AXI_SLAVE_REG[0] <= 32'b0001_00_0000_00_0_1_01_010; //LOADA Row1
        AXI_SLAVE_REG[1] <= 32'b10001_00_0000_01_0_0_01_011; //LOADB Col1
        AXI_SLAVE_REG[2] <= 32'b10101_01_0000_01_0_0_01_011; //LOADB Col2
        AXI_SLAVE_REG[3] <= 32'b11001_10_0000_01_0_0_01_011; //LOADB Col3
        AXI_SLAVE_REG[4] <= 32'b11101_11_0000_01_0_0_01_011; //LOADB Col4
        AXI_SLAVE_REG[5] <= 32'b0000_00_0000_01_0_0_01_100; //MULTACC
        AXI_SLAVE_REG[6] <= 32'b100001_00_0000_00_0_0_01_101; //STORE Row1
        AXI_SLAVE_REG[7] <= 32'b0101_00_0000_00_0_1_01_010; //LOADA Row2
        AXI_SLAVE_REG[8] <= 32'b0000_00_0000_00_0_0_01_100; //MULTACC
        AXI_SLAVE_REG[9] <= 32'b100101_00_0000_00_0_0_01_101; //STORE Row2
        AXI_SLAVE_REG[10] <= 32'b1001_00_0000_00_0_1_01_010; //LOADA Row3
        AXI_SLAVE_REG[11] <= 32'b0000_00_0000_00_0_0_01_100; //MULTACC
        AXI_SLAVE_REG[12] <= 32'b101001_00_0000_00_0_0_01_101; //STORE Row3
        AXI_SLAVE_REG[13] <= 32'b1101_00_0000_00_0_1_01_010; //LOADA Row4
        AXI_SLAVE_REG[14] <= 32'b0000_00_0000_00_0_0_01_100; //MULTACC
        AXI_SLAVE_REG[15] <= 32'b101101_00_0000_00_0_0_01_101; //STORE Row4
        AXI_SLAVE_REG[16] <= 32'b0001_00_0000_00_0_0_00_110; //STOP 
    
        ////////////////////////////////////////////////////////////////////////
        //////////////// 2x2 Matrix Multiplication Instructions ////////////////
        ////////////////////////////////////////////////////////////////////////
 /*   
        AXI_SLAVE_REG[0] <= 32'b0001010001100000010;
        AXI_SLAVE_REG[1] <= 32'b0011000011100000010;
        AXI_SLAVE_REG[2] <= 32'b0101010101110000011;
        AXI_SLAVE_REG[3] <= 32'b0111000111110000011;
        AXI_SLAVE_REG[4] <= 32'b0000000000000000100;
        AXI_SLAVE_REG[5] <= 32'b1001001001000000101;
        AXI_SLAVE_REG[6] <= 32'b0000000000000000110;
        AXI_SLAVE_REG[7] <= 32'b0;
        AXI_SLAVE_REG[8] <= 32'b0;
        AXI_SLAVE_REG[9] <= 32'b0;
        AXI_SLAVE_REG[10] <= 32'b0;
        AXI_SLAVE_REG[11] <= 32'b0;
        AXI_SLAVE_REG[12] <= 32'b0;
        AXI_SLAVE_REG[13] <= 32'b0;
        AXI_SLAVE_REG[14] <= 32'b0;
        AXI_SLAVE_REG[15] <= 32'b0;
        AXI_SLAVE_REG[16] <= 32'b0; */
    end


    assign INSTR_AXI = AXI_SLAVE_REG[PC_AXI];

endmodule