`timescale 1ns/1ps

module Top_PL(
    input logic CLK, RSTN,
    

);


    
endmodule